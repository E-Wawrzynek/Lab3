module OL(
    input [2:0] CurrentState,
    input [1:0] SW,
    input turn_side,
    output [7:0] HEX0,
    output [2:0] LEDR_L,
    output [2:0] LEDR_R
);


endmodule